library verilog;
use verilog.vl_types.all;
entity MIPS_System_tb is
end MIPS_System_tb;
